@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
93 00 00 00 13 01 00 00 93 01 00 00 13 02 00 00
93 02 00 00 13 03 00 00 93 03 00 00 13 04 00 00
93 04 00 00 13 05 00 00 93 05 00 00 13 06 00 00
93 06 00 00 13 07 00 00 93 07 00 00 13 08 00 00
93 08 00 00 13 09 00 00 93 09 00 00 13 0A 00 00
93 0A 00 00 13 0B 00 00 93 0B 00 00 13 0C 00 00
93 0C 00 00 13 0D 00 00 93 0D 00 00 13 0E 00 00
93 0E 00 00 13 0F 00 00 93 0F 00 00 93 00 10 00
13 01 20 00 93 01 30 00 13 02 40 00 93 02 50 00
13 03 60 00 93 03 70 00 13 04 80 00 B3 54 11 40
33 05 64 40 93 55 22 40 13 D6 12 00 93 16 11 00
13 F7 42 00 93 C7 51 00 13 E8 60 00 93 B8 21 00
13 29 52 00 B7 1F 00 00 23 A0 1F 00 23 A2 2F 00
23 A4 3F 00 23 A6 4F 00 23 A8 5F 00 23 AA 6F 00
23 AC 7F 00 23 AE 8F 00 23 A0 9F 02 23 A2 AF 02
23 A4 BF 02 23 A6 CF 02 23 A8 DF 02 23 AA EF 02
23 AC FF 02 23 AE 0F 03 23 A0 1F 05 23 A2 2F 05
83 A8 0F 02 03 A9 4F 02 83 A9 8F 02 03 AA CF 02
83 AA 0F 03 03 AB 4F 03 83 AB 8F 03 03 AC CF 03
83 AC 0F 04 03 AD 4F 04 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 73 00 10 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00
