@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
B7 1F 00 00 93 00 50 00 13 01 A0 00 93 01 B0 FF
13 02 60 FF
