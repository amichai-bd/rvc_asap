@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
93 00 00 00 13 01 00 00 93 01 00 00 13 02 00 00
93 02 00 00 13 03 00 00 93 03 00 00 13 04 00 00
93 04 00 00 13 05 00 00 93 05 00 00 13 06 00 00
93 06 00 00 13 07 00 00 93 07 00 00 13 08 00 00
93 08 00 00 13 09 00 00 93 09 00 00 13 0A 00 00
93 0A 00 00 13 0B 00 00 93 0B 00 00 13 0C 00 00
93 0C 00 00 13 0D 00 00 93 0D 00 00 13 0E 00 00
93 0E 00 00 13 0F 00 00 93 0F 00 00 B7 00 FB FA
93 80 A0 AF 37 C1 BC BC 13 01 C1 CB 93 01 00 00
13 02 00 00 93 02 00 00 13 03 00 00 93 03 00 00
B7 1F 00 00 23 A0 1F 00 23 92 1F 00 23 84 1F 00
23 90 2F 00 83 91 0F 00 03 82 0F 00 83 D2 0F 00
03 C3 0F 00 B7 F3 FA FA 83 A8 0F 02 03 A9 4F 02
83 A9 8F 02 03 AA CF 02 83 AA 0F 03 03 AB 4F 03
83 AB 8F 03 03 AC CF 03 83 AC 0F 04 03 AD 4F 04
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
73 00 10 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00
