@00001000
50 00 00 00 C8 00 00 00 3C 00 00 00 2C 01 00 00
64 00 00 00 46 00 00 00 5A 00 00 00
