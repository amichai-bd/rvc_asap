@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
93 00 00 00 13 01 00 00 93 01 00 00 13 02 00 00
93 02 00 00 13 03 00 00 93 03 00 00 13 04 00 00
93 04 00 00 13 05 00 00 93 05 00 00 13 06 00 00
93 06 00 00 13 07 00 00 93 07 00 00 13 08 00 00
93 08 00 00 13 09 00 00 93 09 00 00 13 0A 00 00
93 0A 00 00 13 0B 00 00 93 0B 00 00 13 0C 00 00
93 0C 00 00 13 0D 00 00 93 0D 00 00 13 0E 00 00
93 0E 00 00 13 0F 00 00 93 0F 00 00 B7 1F 00 00
13 0F 10 00 93 0E 00 00 93 00 10 00 13 01 10 00
93 01 20 00 63 86 20 00 23 A0 DF 01 6F 0E 80 00
23 A0 EF 01 63 96 20 00 23 A2 EF 01 6F 0E 80 00
23 A2 DF 01 63 C6 30 00 23 A4 DF 01 6F 0E 80 00
23 A4 EF 01 63 D6 20 00 23 A6 DF 01 6F 0E 80 00
23 A6 EF 01 63 E6 30 00 23 A8 DF 01 6F 0E 80 00
23 A8 EF 01 63 F6 20 00 23 AA DF 01 6F 0E 80 00
23 AA EF 01 17 F2 FF FF 23 AC 4F 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 73 00 10 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
