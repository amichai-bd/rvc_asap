@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 37 21 00 00
13 01 01 E0 93 81 00 00 13 82 00 00 93 82 00 00
13 83 00 00 93 83 00 00 13 84 00 00 93 84 00 00
13 85 00 00 93 85 00 00 13 86 00 00 93 86 00 00
13 87 00 00 93 87 00 00 13 88 00 00 93 88 00 00
13 89 00 00 93 89 00 00 13 8A 00 00 93 8A 00 00
13 8B 00 00 93 8B 00 00 13 8C 00 00 93 8C 00 00
13 8D 00 00 93 8D 00 00 13 8E 00 00 93 8E 00 00
13 8F 00 00 93 8F 00 00 EF 00 80 00 73 00 10 00
@000000A0
13 01 01 FD 23 26 11 02 23 24 81 02 23 22 91 02
13 04 01 03 B7 17 00 00 93 87 07 00 03 A8 07 00
03 A5 47 00 83 A5 87 00 03 A6 C7 00 83 A6 07 01
03 A7 47 01 83 A7 87 01 23 28 04 FD 23 2A A4 FC
23 2C B4 FC 23 2E C4 FC 23 20 D4 FE 23 22 E4 FE
23 24 F4 FE 93 07 04 FD 93 05 70 00 13 85 07 00
EF 00 80 1B 23 26 04 FE 6F 00 80 03 83 27 C4 FE
13 97 27 00 B7 17 00 00 33 07 F7 00 83 27 C4 FE
93 97 27 00 93 06 04 FF B3 87 F6 00 83 A7 07 FE
23 20 F7 00 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 C4 FE 93 07 60 00 E3 D2 E7 FC B7 17 00 00
93 84 C7 01 13 05 90 00 EF 00 40 0A 93 07 05 00
23 A0 F4 00 B7 17 00 00 93 84 07 02 93 05 00 01
13 05 80 01 EF 00 80 02 93 07 05 00 23 A0 F4 00
93 07 00 00 13 85 07 00 83 20 C1 02 03 24 81 02
83 24 41 02 13 01 01 03 67 80 00 00 13 01 01 FE
23 2E 11 00 23 2C 81 00 13 04 01 02 23 26 A4 FE
23 24 B4 FE 83 27 84 FE 63 86 07 02 83 27 C4 FE
83 25 84 FE 13 85 07 00 EF 00 40 25 93 07 05 00
93 85 07 00 03 25 84 FE EF F0 5F FC 93 07 05 00
6F 00 80 00 83 27 C4 FE 13 85 07 00 83 20 C1 01
03 24 81 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 11 00 23 2C 81 00 23 2A 91 00 13 04 01 02
23 26 A4 FE 03 27 C4 FE 93 07 10 00 63 E6 E7 00
83 27 C4 FE 6F 00 00 03 83 27 C4 FE 93 87 F7 FF
13 85 07 00 EF F0 9F FC 93 04 05 00 83 27 C4 FE
93 87 E7 FF 13 85 07 00 EF F0 5F FB 93 07 05 00
B3 87 F4 00 13 85 07 00 83 20 C1 01 03 24 81 01
83 24 41 01 13 01 01 02 67 80 00 00 13 01 01 FD
23 26 81 02 13 04 01 03 23 2E A4 FC 23 2C B4 FC
83 27 C4 FD 83 A7 07 00 23 26 F4 FE 83 27 84 FD
03 A7 07 00 83 27 C4 FD 23 A0 E7 00 83 27 84 FD
03 27 C4 FE 23 A0 E7 00 13 00 00 00 03 24 C1 02
13 01 01 03 67 80 00 00 13 01 01 FD 23 26 11 02
23 24 81 02 13 04 01 03 23 2E A4 FC 23 2C B4 FC
23 26 04 FE 6F 00 C0 09 23 24 04 FE 6F 00 00 07
83 27 84 FE 93 97 27 00 03 27 C4 FD B3 07 F7 00
03 A7 07 00 83 27 84 FE 93 87 17 00 93 97 27 00
83 26 C4 FD B3 87 F6 00 83 A7 07 00 63 DA E7 02
83 27 84 FE 93 97 27 00 03 27 C4 FD B3 06 F7 00
83 27 84 FE 93 87 17 00 93 97 27 00 03 27 C4 FD
B3 07 F7 00 93 85 07 00 13 85 06 00 EF F0 1F F3
83 27 84 FE 93 87 17 00 23 24 F4 FE 03 27 84 FD
83 27 C4 FE B3 07 F7 40 93 87 F7 FF 03 27 84 FE
E3 40 F7 F8 83 27 C4 FE 93 87 17 00 23 26 F4 FE
83 27 84 FD 93 87 F7 FF 03 27 C4 FE E3 4E F7 F4
13 00 00 00 13 00 00 00 83 20 C1 02 03 24 81 02
13 01 01 03 67 80 00 00 63 40 05 06 63 C6 05 06
13 86 05 00 93 05 05 00 13 05 F0 FF 63 0C 06 02
93 06 10 00 63 7A B6 00 63 58 C0 00 13 16 16 00
93 96 16 00 E3 6A B6 FE 13 05 00 00 63 E6 C5 00
B3 85 C5 40 33 65 D5 00 93 D6 16 00 13 56 16 00
E3 96 06 FE 67 80 00 00 93 82 00 00 EF F0 5F FB
13 85 05 00 67 80 02 00 33 05 A0 40 63 48 B0 00
B3 05 B0 40 6F F0 DF F9 B3 05 B0 40 93 82 00 00
EF F0 1F F9 33 05 A0 40 67 80 02 00 93 82 00 00
63 CA 05 00 63 4C 05 00 EF F0 9F F7 13 85 05 00
67 80 02 00 B3 05 B0 40 E3 58 05 FE 33 05 A0 40
EF F0 1F F6 33 05 B0 40 67 80 02 00
