module test (
    input  logic in_0,
    input  logic in_1,
    output logic out
);
assign out = in_0 & in_1;
endmodule