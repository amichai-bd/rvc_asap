@00001000
01 00 00 00 02 00 00 00 03 00 00 00 04 00 00 00
