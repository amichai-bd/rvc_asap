@00001000
