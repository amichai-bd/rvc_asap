@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 37 21 00 00
13 01 01 E0 93 81 00 00 13 82 00 00 93 82 00 00
13 83 00 00 93 83 00 00 13 84 00 00 93 84 00 00
13 85 00 00 93 85 00 00 13 86 00 00 93 86 00 00
13 87 00 00 93 87 00 00 13 88 00 00 93 88 00 00
13 89 00 00 93 89 00 00 13 8A 00 00 93 8A 00 00
13 8B 00 00 93 8B 00 00 13 8C 00 00 93 8C 00 00
13 8D 00 00 93 8D 00 00 13 8E 00 00 93 8E 00 00
13 8F 00 00 93 8F 00 00 EF 00 80 03 73 00 10 00
@000000A0
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 A4 FE
23 24 B4 FE 03 27 C4 FE 83 27 84 FE B3 07 F7 00
13 85 07 00 03 24 C1 01 13 01 01 02 67 80 00 00
13 01 01 FD 23 26 11 02 23 24 81 02 13 04 01 03
B7 17 00 00 93 87 07 00 03 A6 07 00 83 A6 47 00
03 A7 87 00 83 A7 C7 00 23 2A C4 FC 23 2C D4 FC
23 2E E4 FC 23 20 F4 FE 93 07 30 00 23 26 F4 FE
93 07 50 00 23 24 F4 FE 83 25 84 FE 03 25 C4 FE
EF F0 1F F8 23 22 A4 FE 93 07 00 00 13 85 07 00
83 20 C1 02 03 24 81 02 13 01 01 03 67 80 00 00
