@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 37 21 00 00 EF 00 40 04 73 00 10 00
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 23 26 04 FE 03 27 C4 FD 83 27 84 FD
B3 07 F7 00 23 26 F4 FE 83 27 C4 FE 13 85 07 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FE
23 2E 11 00 23 2C 81 00 13 04 01 02 93 07 20 00
23 26 F4 FE 93 07 40 00 23 24 F4 FE 83 25 84 FE
03 25 C4 FE EF F0 DF F9 23 22 A4 FE 93 07 00 00
13 85 07 00 83 20 C1 01 03 24 81 01 13 01 01 02
67 80 00 00
